----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/27/2024 11:45:36 PM
-- Design Name: 
-- Module Name: hdmi_pixel_pusher - hdmi_pixel_pusher_arch
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity hdmi_pixel_pusher is
    Port ( clk, clk_en, VS : in STD_LOGIC := '0';
         pixel : in STD_LOGIC_VECTOR (7 downto 0);
         hcount : in STD_LOGIC_VECTOR (9 downto 0) := (others => '0');
         vid : in STD_LOGIC := '0';
         R, B : out STD_LOGIC_VECTOR (4 downto 0) := (others => '0');
         G : out STD_LOGIC_VECTOR (5 downto 0) := (others => '0');
         addr : out STD_LOGIC_VECTOR (17 downto 0);
         hdmiOut : out std_logic_vector(23 downto 0));
end hdmi_pixel_pusher;

architecture hdmi_pixel_pusher_arch of hdmi_pixel_pusher is

    signal addr_Reg : std_logic_vector(17 downto 0);
    signal red, blue : std_logic_vector(4 downto 0);
    signal green : std_logic_vector(5 downto 0);
begin

    addr <= addr_Reg;

    hdmiOut <= Red & "000" & Blue & "000" & Green & "00";
    addr_proc : process(clk) begin
        if(rising_edge(clk)) then
            if(VS = '0') then
                addr_Reg  <= (others => '0');
            end if;
            if(clk_en = '1' and vid = '1' and unsigned(hcount)<480) then
                addr_Reg <= std_logic_vector(unsigned(addr_Reg)+1);
                R <= pixel(7 downto 5) & "00";
                G <= pixel(4 downto 2) & "000";
                B <= pixel(1 downto 0) & "000";
                Red <= pixel(7 downto 5) & "00";
                Green <= pixel(4 downto 2) & "000";
                Blue <= pixel(1 downto 0) & "000";
            elsif(clk_en = '1' and vid = '1' and unsigned(hcount)>=480) then
                R <= (others => '0');
                B <= (others => '0');
                G <= (others => '0');
                Red <= (others => '0');
                Blue <= (others => '0');
                Green <= (others => '0');
            end if;
        end if;
    end process addr_proc;
end hdmi_pixel_pusher_arch;